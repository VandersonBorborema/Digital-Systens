library verilog;
use verilog.vl_types.all;
entity processador16bits_vlg_vec_tst is
end processador16bits_vlg_vec_tst;
