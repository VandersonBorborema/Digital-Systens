library verilog;
use verilog.vl_types.all;
entity somador_4bits_vlg_vec_tst is
end somador_4bits_vlg_vec_tst;
